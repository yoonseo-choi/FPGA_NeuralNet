module sigmoid (input [15:0] h0,
                output logic out
)